VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO tt_um_collosal_demo
  CLASS BLOCK ;
  FOREIGN tt_um_collosal_demo ;
  ORIGIN 0.000 0.000 ;
  SIZE 856.520 BY 511.360 ;
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 21.580 2.480 23.180 508.880 ;
    END
    PORT
      LAYER met4 ;
        RECT 60.450 2.480 62.050 508.880 ;
    END
    PORT
      LAYER met4 ;
        RECT 99.320 2.480 100.920 508.880 ;
    END
    PORT
      LAYER met4 ;
        RECT 138.190 2.480 139.790 508.880 ;
    END
    PORT
      LAYER met4 ;
        RECT 177.060 2.480 178.660 508.880 ;
    END
    PORT
      LAYER met4 ;
        RECT 215.930 2.480 217.530 508.880 ;
    END
    PORT
      LAYER met4 ;
        RECT 254.800 2.480 256.400 508.880 ;
    END
    PORT
      LAYER met4 ;
        RECT 293.670 2.480 295.270 508.880 ;
    END
    PORT
      LAYER met4 ;
        RECT 332.540 2.480 334.140 508.880 ;
    END
    PORT
      LAYER met4 ;
        RECT 371.410 2.480 373.010 508.880 ;
    END
    PORT
      LAYER met4 ;
        RECT 410.280 2.480 411.880 508.880 ;
    END
    PORT
      LAYER met4 ;
        RECT 449.150 2.480 450.750 508.880 ;
    END
    PORT
      LAYER met4 ;
        RECT 488.020 2.480 489.620 508.880 ;
    END
    PORT
      LAYER met4 ;
        RECT 526.890 2.480 528.490 508.880 ;
    END
    PORT
      LAYER met4 ;
        RECT 565.760 2.480 567.360 508.880 ;
    END
    PORT
      LAYER met4 ;
        RECT 604.630 2.480 606.230 508.880 ;
    END
    PORT
      LAYER met4 ;
        RECT 643.500 2.480 645.100 508.880 ;
    END
    PORT
      LAYER met4 ;
        RECT 682.370 2.480 683.970 508.880 ;
    END
    PORT
      LAYER met4 ;
        RECT 721.240 2.480 722.840 508.880 ;
    END
    PORT
      LAYER met4 ;
        RECT 760.110 2.480 761.710 508.880 ;
    END
    PORT
      LAYER met4 ;
        RECT 798.980 2.480 800.580 508.880 ;
    END
    PORT
      LAYER met4 ;
        RECT 837.850 2.480 839.450 508.880 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 18.280 2.480 19.880 508.880 ;
    END
    PORT
      LAYER met4 ;
        RECT 57.150 2.480 58.750 508.880 ;
    END
    PORT
      LAYER met4 ;
        RECT 96.020 2.480 97.620 508.880 ;
    END
    PORT
      LAYER met4 ;
        RECT 134.890 2.480 136.490 508.880 ;
    END
    PORT
      LAYER met4 ;
        RECT 173.760 2.480 175.360 508.880 ;
    END
    PORT
      LAYER met4 ;
        RECT 212.630 2.480 214.230 508.880 ;
    END
    PORT
      LAYER met4 ;
        RECT 251.500 2.480 253.100 508.880 ;
    END
    PORT
      LAYER met4 ;
        RECT 290.370 2.480 291.970 508.880 ;
    END
    PORT
      LAYER met4 ;
        RECT 329.240 2.480 330.840 508.880 ;
    END
    PORT
      LAYER met4 ;
        RECT 368.110 2.480 369.710 508.880 ;
    END
    PORT
      LAYER met4 ;
        RECT 406.980 2.480 408.580 508.880 ;
    END
    PORT
      LAYER met4 ;
        RECT 445.850 2.480 447.450 508.880 ;
    END
    PORT
      LAYER met4 ;
        RECT 484.720 2.480 486.320 508.880 ;
    END
    PORT
      LAYER met4 ;
        RECT 523.590 2.480 525.190 508.880 ;
    END
    PORT
      LAYER met4 ;
        RECT 562.460 2.480 564.060 508.880 ;
    END
    PORT
      LAYER met4 ;
        RECT 601.330 2.480 602.930 508.880 ;
    END
    PORT
      LAYER met4 ;
        RECT 640.200 2.480 641.800 508.880 ;
    END
    PORT
      LAYER met4 ;
        RECT 679.070 2.480 680.670 508.880 ;
    END
    PORT
      LAYER met4 ;
        RECT 717.940 2.480 719.540 508.880 ;
    END
    PORT
      LAYER met4 ;
        RECT 756.810 2.480 758.410 508.880 ;
    END
    PORT
      LAYER met4 ;
        RECT 795.680 2.480 797.280 508.880 ;
    END
    PORT
      LAYER met4 ;
        RECT 834.550 2.480 836.150 508.880 ;
    END
  END VPWR
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 143.830 510.360 144.130 511.360 ;
    END
  END clk
  PIN ena
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 146.590 510.360 146.890 511.360 ;
    END
  END ena
  PIN rst_n
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met4 ;
        RECT 141.070 510.360 141.370 511.360 ;
    END
  END rst_n
  PIN ui_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met4 ;
        RECT 138.310 510.360 138.610 511.360 ;
    END
  END ui_in[0]
  PIN ui_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met4 ;
        RECT 135.550 510.360 135.850 511.360 ;
    END
  END ui_in[1]
  PIN ui_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met4 ;
        RECT 132.790 510.360 133.090 511.360 ;
    END
  END ui_in[2]
  PIN ui_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met4 ;
        RECT 130.030 510.360 130.330 511.360 ;
    END
  END ui_in[3]
  PIN ui_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 127.270 510.360 127.570 511.360 ;
    END
  END ui_in[4]
  PIN ui_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 124.510 510.360 124.810 511.360 ;
    END
  END ui_in[5]
  PIN ui_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met4 ;
        RECT 121.750 510.360 122.050 511.360 ;
    END
  END ui_in[6]
  PIN ui_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 118.990 510.360 119.290 511.360 ;
    END
  END ui_in[7]
  PIN uio_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met4 ;
        RECT 116.230 510.360 116.530 511.360 ;
    END
  END uio_in[0]
  PIN uio_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met4 ;
        RECT 113.470 510.360 113.770 511.360 ;
    END
  END uio_in[1]
  PIN uio_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met4 ;
        RECT 110.710 510.360 111.010 511.360 ;
    END
  END uio_in[2]
  PIN uio_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 107.950 510.360 108.250 511.360 ;
    END
  END uio_in[3]
  PIN uio_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met4 ;
        RECT 105.190 510.360 105.490 511.360 ;
    END
  END uio_in[4]
  PIN uio_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met4 ;
        RECT 102.430 510.360 102.730 511.360 ;
    END
  END uio_in[5]
  PIN uio_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met4 ;
        RECT 99.670 510.360 99.970 511.360 ;
    END
  END uio_in[6]
  PIN uio_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met4 ;
        RECT 96.910 510.360 97.210 511.360 ;
    END
  END uio_in[7]
  PIN uio_oe[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met4 ;
        RECT 49.990 510.360 50.290 511.360 ;
    END
  END uio_oe[0]
  PIN uio_oe[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met4 ;
        RECT 47.230 510.360 47.530 511.360 ;
    END
  END uio_oe[1]
  PIN uio_oe[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met4 ;
        RECT 44.470 510.360 44.770 511.360 ;
    END
  END uio_oe[2]
  PIN uio_oe[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met4 ;
        RECT 41.710 510.360 42.010 511.360 ;
    END
  END uio_oe[3]
  PIN uio_oe[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met4 ;
        RECT 38.950 510.360 39.250 511.360 ;
    END
  END uio_oe[4]
  PIN uio_oe[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met4 ;
        RECT 36.190 510.360 36.490 511.360 ;
    END
  END uio_oe[5]
  PIN uio_oe[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met4 ;
        RECT 33.430 510.360 33.730 511.360 ;
    END
  END uio_oe[6]
  PIN uio_oe[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met4 ;
        RECT 30.670 510.360 30.970 511.360 ;
    END
  END uio_oe[7]
  PIN uio_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met4 ;
        RECT 72.070 510.360 72.370 511.360 ;
    END
  END uio_out[0]
  PIN uio_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met4 ;
        RECT 69.310 510.360 69.610 511.360 ;
    END
  END uio_out[1]
  PIN uio_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met4 ;
        RECT 66.550 510.360 66.850 511.360 ;
    END
  END uio_out[2]
  PIN uio_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met4 ;
        RECT 63.790 510.360 64.090 511.360 ;
    END
  END uio_out[3]
  PIN uio_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met4 ;
        RECT 61.030 510.360 61.330 511.360 ;
    END
  END uio_out[4]
  PIN uio_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met4 ;
        RECT 58.270 510.360 58.570 511.360 ;
    END
  END uio_out[5]
  PIN uio_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met4 ;
        RECT 55.510 510.360 55.810 511.360 ;
    END
  END uio_out[6]
  PIN uio_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met4 ;
        RECT 52.750 510.360 53.050 511.360 ;
    END
  END uio_out[7]
  PIN uo_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met4 ;
        RECT 94.150 510.360 94.450 511.360 ;
    END
  END uo_out[0]
  PIN uo_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met4 ;
        RECT 91.390 510.360 91.690 511.360 ;
    END
  END uo_out[1]
  PIN uo_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met4 ;
        RECT 88.630 510.360 88.930 511.360 ;
    END
  END uo_out[2]
  PIN uo_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met4 ;
        RECT 85.870 510.360 86.170 511.360 ;
    END
  END uo_out[3]
  PIN uo_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met4 ;
        RECT 83.110 510.360 83.410 511.360 ;
    END
  END uo_out[4]
  PIN uo_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met4 ;
        RECT 80.350 510.360 80.650 511.360 ;
    END
  END uo_out[5]
  PIN uo_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met4 ;
        RECT 77.590 510.360 77.890 511.360 ;
    END
  END uo_out[6]
  PIN uo_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met4 ;
        RECT 74.830 510.360 75.130 511.360 ;
    END
  END uo_out[7]
  OBS
      LAYER li1 ;
        RECT 2.760 2.635 853.760 508.725 ;
      LAYER met1 ;
        RECT 2.460 2.080 854.060 510.980 ;
      LAYER met2 ;
        RECT 4.240 2.050 853.200 511.010 ;
      LAYER met3 ;
        RECT 11.105 2.555 851.855 510.505 ;
      LAYER met4 ;
        RECT 31.370 509.960 33.030 511.010 ;
        RECT 34.130 509.960 35.790 511.010 ;
        RECT 36.890 509.960 38.550 511.010 ;
        RECT 39.650 509.960 41.310 511.010 ;
        RECT 42.410 509.960 44.070 511.010 ;
        RECT 45.170 509.960 46.830 511.010 ;
        RECT 47.930 509.960 49.590 511.010 ;
        RECT 50.690 509.960 52.350 511.010 ;
        RECT 53.450 509.960 55.110 511.010 ;
        RECT 56.210 509.960 57.870 511.010 ;
        RECT 58.970 509.960 60.630 511.010 ;
        RECT 61.730 509.960 63.390 511.010 ;
        RECT 64.490 509.960 66.150 511.010 ;
        RECT 67.250 509.960 68.910 511.010 ;
        RECT 70.010 509.960 71.670 511.010 ;
        RECT 72.770 509.960 74.430 511.010 ;
        RECT 75.530 509.960 77.190 511.010 ;
        RECT 78.290 509.960 79.950 511.010 ;
        RECT 81.050 509.960 82.710 511.010 ;
        RECT 83.810 509.960 85.470 511.010 ;
        RECT 86.570 509.960 88.230 511.010 ;
        RECT 89.330 509.960 90.990 511.010 ;
        RECT 92.090 509.960 93.750 511.010 ;
        RECT 94.850 509.960 96.510 511.010 ;
        RECT 97.610 509.960 99.270 511.010 ;
        RECT 100.370 509.960 102.030 511.010 ;
        RECT 103.130 509.960 104.790 511.010 ;
        RECT 105.890 509.960 107.550 511.010 ;
        RECT 108.650 509.960 110.310 511.010 ;
        RECT 111.410 509.960 113.070 511.010 ;
        RECT 114.170 509.960 115.830 511.010 ;
        RECT 116.930 509.960 118.590 511.010 ;
        RECT 119.690 509.960 121.350 511.010 ;
        RECT 122.450 509.960 124.110 511.010 ;
        RECT 125.210 509.960 126.870 511.010 ;
        RECT 127.970 509.960 129.630 511.010 ;
        RECT 130.730 509.960 132.390 511.010 ;
        RECT 133.490 509.960 135.150 511.010 ;
        RECT 136.250 509.960 137.910 511.010 ;
        RECT 139.010 509.960 140.670 511.010 ;
        RECT 141.770 509.960 143.430 511.010 ;
        RECT 144.530 509.960 146.190 511.010 ;
        RECT 147.290 509.960 806.545 511.010 ;
        RECT 30.655 509.280 806.545 509.960 ;
        RECT 30.655 15.135 56.750 509.280 ;
        RECT 59.150 15.135 60.050 509.280 ;
        RECT 62.450 15.135 95.620 509.280 ;
        RECT 98.020 15.135 98.920 509.280 ;
        RECT 101.320 15.135 134.490 509.280 ;
        RECT 136.890 15.135 137.790 509.280 ;
        RECT 140.190 15.135 173.360 509.280 ;
        RECT 175.760 15.135 176.660 509.280 ;
        RECT 179.060 15.135 212.230 509.280 ;
        RECT 214.630 15.135 215.530 509.280 ;
        RECT 217.930 15.135 251.100 509.280 ;
        RECT 253.500 15.135 254.400 509.280 ;
        RECT 256.800 15.135 289.970 509.280 ;
        RECT 292.370 15.135 293.270 509.280 ;
        RECT 295.670 15.135 328.840 509.280 ;
        RECT 331.240 15.135 332.140 509.280 ;
        RECT 334.540 15.135 367.710 509.280 ;
        RECT 370.110 15.135 371.010 509.280 ;
        RECT 373.410 15.135 406.580 509.280 ;
        RECT 408.980 15.135 409.880 509.280 ;
        RECT 412.280 15.135 445.450 509.280 ;
        RECT 447.850 15.135 448.750 509.280 ;
        RECT 451.150 15.135 484.320 509.280 ;
        RECT 486.720 15.135 487.620 509.280 ;
        RECT 490.020 15.135 523.190 509.280 ;
        RECT 525.590 15.135 526.490 509.280 ;
        RECT 528.890 15.135 562.060 509.280 ;
        RECT 564.460 15.135 565.360 509.280 ;
        RECT 567.760 15.135 600.930 509.280 ;
        RECT 603.330 15.135 604.230 509.280 ;
        RECT 606.630 15.135 639.800 509.280 ;
        RECT 642.200 15.135 643.100 509.280 ;
        RECT 645.500 15.135 678.670 509.280 ;
        RECT 681.070 15.135 681.970 509.280 ;
        RECT 684.370 15.135 717.540 509.280 ;
        RECT 719.940 15.135 720.840 509.280 ;
        RECT 723.240 15.135 756.410 509.280 ;
        RECT 758.810 15.135 759.710 509.280 ;
        RECT 762.110 15.135 795.280 509.280 ;
        RECT 797.680 15.135 798.580 509.280 ;
        RECT 800.980 15.135 806.545 509.280 ;
  END
END tt_um_collosal_demo
END LIBRARY

